netcdf sample {
dimensions:
	lon = 10 ;
	lat = 10 ;
	count = 10 ;
	city = 10 ;
	time = UNLIMITED ; // (10 currently)
variables:
	float Longitude(lon) ;
	float Latitude(lat) ;
	int Time(time) ;
	string City(city) ;
	int wikipediaWC(count) ;
	float population(time, lon, lat) ;
	float populationCity(time, city) ;
data:

 Longitude = 90.48157, 89.69103, 63.87073, 82.37345, 77.51483, 74.39978, 
    59.75166, 73.70914, 57.59724, 92.57875 ;

 Latitude = 6.505907, -19.88314, -2.398372, 18.44205, 21.24537, -22.44801, 
    -24.80032, 11.25267, 17.59253, -1.663467 ;

 Time = 737463, 737303, 737151, 737265, 737857, 737539, 737124, 737426, 
    737718, 736869 ;

 City = "Amsterdam", "Barcelona", "Paris", "Geneva", "Munich", "Athens", 
    "Vienna", "Karachi", "Islamabad", "Multan" ;

 wikipediaWC = 70, 1, 86, 34, 24, 5, 23, 85, 71, 73 ;

 population =
  2861476, 4796172, 3939779, 2174007, 1524640, 1703603, 3007837, 2827959, 
    279045, 703039,
  476287, 4624334, 2338709, 2001613, 3676067, 218482, 2956042, 4684129, 
    1968832, 2468503,
  1108385, 2359834, 4348155, 1950685, 2928051, 4759547, 1649550, 1375366, 
    4812150, 2962571,
  2209303, 2425839, 3364742, 313462, 1631201, 1285396, 4968936, 2613729, 
    993485, 2420379,
  728479, 4616190, 1248444, 3073380, 4793090, 1516225, 4518731, 1967001, 
    1900529, 961992,
  1980208, 2964583, 1527357, 3785738, 1402342, 4022199, 970944, 3254604, 
    1147930, 3656873,
  3071387, 408691, 538235, 3017468, 2895795, 564453, 1460631, 2553834, 
    4747282, 798694,
  4706551, 2159667, 1785089, 4514280, 3760451, 521993, 3893586, 3275774, 
    1890205, 2565699,
  3981712, 4178629, 355623, 2255359, 1599420, 2929999, 1073225, 1436748, 
    3407535, 4536919,
  67241, 4517967, 812780, 512066, 3290481, 1807625, 2535234, 3084976, 660646, 
    3123796,
  2835446, 1493169, 348551, 3407874, 4202085, 2434216, 1861140, 4909047, 
    1132778, 3240212,
  1333470, 1053196, 263334, 437085, 3523291, 4119038, 3418270, 3665349, 
    1860651, 3151399,
  238162, 4154454, 2385030, 1604966, 1428613, 879374, 2132691, 4880438, 
    3761556, 4641167,
  1879566, 2997716, 715376, 3756578, 1770880, 559445, 2378974, 2632380, 
    3000405, 702681,
  459343, 4771769, 1795472, 4507013, 4352325, 2553857, 197061, 110172, 
    1451632, 2643427,
  1170791, 3192446, 857804, 339909, 262709, 619882, 4931912, 1953899, 
    4461786, 2923550,
  4452465, 316792, 3567531, 3050143, 3996072, 315351, 345214, 4938606, 
    2718115, 4596810,
  4465670, 3286750, 3936053, 2431468, 540160, 1020748, 2356166, 4132852, 
    1226967, 3167523,
  1283299, 3645368, 3306941, 2838591, 964917, 2145977, 2214226, 2693514, 
    3180774, 699573,
  1377860, 255655, 1938112, 2819024, 3846825, 1623224, 2808310, 4224494, 
    929362, 2017191,
  4009053, 4926510, 2098719, 2778439, 3493972, 3297482, 1681269, 2630725, 
    4742822, 315366,
  4411464, 4881162, 470724, 447949, 4830835, 2655159, 4964896, 4320586, 
    3893803, 3916602,
  3704721, 794659, 3990744, 3893877, 4214824, 838040, 3978033, 754021, 
    3422378, 60947,
  194199, 1616989, 3269260, 4051893, 133047, 1852259, 1627194, 3877905, 
    3741497, 4979135,
  2320162, 946236, 3342466, 4363474, 2559264, 2550549, 4308859, 795641, 
    2524245, 1648404,
  2544177, 1763662, 1865145, 346416, 4631360, 2398686, 1073679, 4968995, 
    1242051, 1376234,
  3050880, 897004, 2898690, 2183829, 4579340, 4571431, 4731620, 3393779, 
    4644356, 2561553,
  1521185, 4259016, 2371033, 196115, 756879, 2559483, 1169720, 4035901, 
    355488, 2539326,
  2187412, 1084733, 2409884, 3174132, 3933430, 3376000, 2931143, 1004463, 
    3953755, 213405,
  2651204, 3763733, 3074157, 2045081, 1901294, 4326903, 2810740, 1300735, 
    2107413, 1504679,
  4288159, 3542186, 4440453, 3484492, 4799193, 1981880, 1021989, 2839647, 
    1174829, 883268,
  2986478, 111392, 3912474, 4300551, 1043676, 2276096, 1589483, 806400, 
    597729, 4919184,
  4970705, 3499209, 341751, 1830933, 3610639, 1430343, 4309507, 4971171, 
    816435, 1801584,
  1454354, 1713956, 2067978, 4955707, 4535492, 3661784, 3352472, 3155814, 
    4456604, 4686606,
  4890553, 3697537, 4943850, 16904, 3925780, 3027856, 1667294, 682378, 
    2238416, 2662444,
  2934885, 1337032, 4706442, 629500, 1818577, 2105469, 885017, 258637, 
    3904684, 2257689,
  1454161, 2572917, 863765, 1876496, 4550242, 3422456, 2248390, 1801236, 
    4412877, 3199452,
  3940583, 2435723, 4385169, 3118375, 1192536, 4857741, 3773779, 3618767, 
    2914579, 3529304,
  3104249, 3934420, 3762305, 1263742, 4857843, 1301547, 1600326, 2293967, 
    4480313, 283142,
  391405, 4786974, 4086708, 362065, 4892758, 1822178, 2695005, 3375974, 
    4542848, 70336,
  3349287, 249326, 1272822, 879515, 64452, 4322136, 432530, 4407113, 4743467, 
    488349,
  2015926, 3964073, 4526284, 227797, 320455, 3573053, 2387004, 3115058, 
    2359621, 4665346,
  2910249, 2768280, 1784270, 4387346, 4149456, 2572901, 2452425, 957922, 
    2630627, 192958,
  3566278, 130883, 1007027, 3899727, 593840, 4074080, 1807234, 923521, 
    3295362, 4186505,
  2769301, 3829348, 1630450, 3860970, 3740387, 150938, 3788904, 3624831, 
    2253704, 2823937,
  2311119, 370419, 707616, 3740540, 3849261, 4523060, 2697497, 539694, 
    3474334, 3608845,
  974335, 147653, 919838, 1241281, 1703885, 1045750, 985446, 2727713, 
    3626393, 2095913,
  43078, 1403201, 544622, 1773476, 3051775, 2441546, 4058259, 2762759, 
    3366189, 3381864,
  2182202, 4421686, 3535886, 2034297, 872420, 521802, 3648964, 2463404, 
    3750172, 852328,
  2965561, 111073, 791049, 2274262, 2398799, 473033, 2474625, 2942114, 
    2566268, 3884208,
  3307683, 4895029, 1678761, 4889720, 4669999, 4456521, 4130847, 4257203, 
    485946, 1660574,
  4275052, 3049396, 4899872, 498124, 3971186, 4729117, 3322129, 1820506, 
    3019439, 644180,
  3383049, 4738238, 673477, 1677922, 4407879, 1528536, 4160772, 3443889, 
    1867849, 1185573,
  259958, 2667373, 1986851, 1148316, 4929862, 3662372, 3250478, 1498557, 
    4554936, 130962,
  2602715, 13467, 3740964, 3897525, 1082318, 2757589, 3526030, 1388978, 
    4861798, 2915625,
  373956, 2097042, 3050945, 3625501, 2598121, 583387, 1322725, 4526418, 
    1508255, 4621545,
  2968745, 3202732, 3158655, 188441, 827255, 2525197, 1478129, 2440348, 
    1965447, 1116428,
  831620, 4780633, 4908636, 3748580, 2909355, 974427, 527758, 3874681, 
    2702692, 1699743,
  172205, 3946661, 4809315, 3319473, 2088906, 677325, 541570, 171834, 912495, 
    4615898,
  2698297, 3042216, 4068266, 531300, 3842055, 2785083, 1894147, 2993947, 
    3445858, 2158669,
  1194060, 3104932, 1547439, 3690805, 4880042, 2350909, 665237, 410079, 
    245691, 697402,
  3969706, 2677074, 3904302, 3328160, 102280, 1078689, 450552, 2483658, 
    1680688, 1350037,
  2556754, 4774327, 2181629, 3229289, 1368292, 1784041, 4089792, 3334537, 
    3681588, 2503518,
  137875, 1166830, 3172661, 541419, 1257366, 3666370, 1214557, 1687943, 
    4867731, 2272011,
  1447321, 1301825, 1070026, 3775533, 3920228, 1005640, 1144331, 1904469, 
    2883123, 3913268,
  754412, 1041399, 1516750, 1658640, 2179861, 3895077, 2117741, 4619658, 
    4966021, 4300177,
  569027, 1748507, 2293821, 3390373, 888435, 2040716, 1303244, 4817072, 
    1237442, 3616985,
  251056, 945584, 1368869, 227459, 744678, 963861, 2238210, 4376764, 572841, 
    1544760,
  1890294, 4930783, 2152613, 4376575, 2429645, 3577175, 3865681, 1662660, 
    944782, 2647375,
  3443178, 4435596, 601330, 15237, 2390178, 3256482, 178146, 4277353, 923063, 
    4909837,
  4974637, 45020, 3507745, 1841481, 861250, 4636488, 1839112, 1150827, 
    3036215, 1717563,
  4479242, 3156304, 1064074, 1599996, 2455095, 263276, 2772011, 410836, 
    2411289, 1199126,
  1341890, 832269, 1275690, 24095, 2476972, 1824677, 4232347, 1979591, 
    2618693, 4008773,
  2755523, 4321157, 4878443, 4832173, 2669567, 2931072, 2112715, 2278911, 
    1896732, 4114952,
  4720470, 4601565, 2931174, 571546, 2719479, 1392854, 4201914, 928464, 
    3934399, 1142970,
  4964128, 720584, 1242547, 287517, 3150268, 4254114, 2791464, 212118, 
    4860427, 4373660,
  1262598, 2895721, 3929475, 4060985, 822857, 4998787, 4024389, 644093, 
    2763386, 1061289,
  2063060, 342221, 1311233, 207880, 1716129, 1361117, 3971263, 1600832, 
    3149236, 2912732,
  4119865, 3112308, 1538108, 4495841, 2592032, 1348672, 2656670, 3553221, 
    385384, 960143,
  3246789, 3196962, 1425860, 4132745, 282668, 4245608, 4158010, 3760370, 
    2597232, 4227287,
  3522717, 845722, 2934883, 2000171, 1242906, 3696928, 1280176, 2341328, 
    848715, 1778339,
  4690416, 2390014, 2268439, 561977, 4826427, 2019185, 1624185, 1361260, 
    356517, 4866860,
  2776344, 3390030, 2642429, 2669721, 3852565, 3033257, 3167419, 1652194, 
    94581, 3637510,
  494463, 4100898, 298828, 1248939, 1361276, 3016404, 1654437, 3468195, 
    4678495, 2393320,
  3963875, 2853511, 3714456, 4439099, 4589708, 2834331, 2720981, 4153494, 
    4891300, 2163110,
  357311, 3892417, 556017, 460917, 1077203, 4929159, 2383307, 695529, 532595, 
    4733213,
  714298, 3560473, 873434, 1219090, 2122550, 4159324, 4244149, 676449, 
    4098811, 2437246,
  2691553, 2715247, 3233409, 159954, 3401422, 3415334, 3103505, 2474154, 
    3416896, 839384,
  2559484, 1954276, 240016, 1640953, 279822, 3142054, 1896166, 3501090, 
    2267987, 2802713,
  1620520, 1016264, 1384185, 3311185, 4147918, 627416, 3912816, 1923431, 
    4755093, 1542830,
  2987042, 563966, 1212285, 3247038, 4172673, 4386152, 1218520, 1771868, 
    3334642, 4856037,
  1112626, 2617595, 3647825, 3875823, 2092709, 3749329, 1759817, 3324275, 
    4259848, 2742739,
  1648302, 3198385, 1207325, 2451122, 2218810, 2544069, 4530387, 804682, 
    1111271, 4605487,
  2663575, 4972473, 4093494, 1009906, 3828682, 766011, 4710288, 4503504, 
    2849103, 3191226,
  274842, 676396, 512619, 4764428, 3735992, 2875656, 583951, 1206257, 
    4371022, 413199,
  4273444, 197999, 851739, 2198683, 4556872, 2362048, 4457861, 760046, 
    3754461, 1787647,
  2834617, 3181762, 3896941, 274279, 2331361, 2953760, 1035689, 2011202, 
    2857722, 3123417,
  2713968, 4002238, 3156947, 2813635, 4310340, 4513590, 4514116, 4085112, 
    2562496, 847127,
  3938828, 3028731, 4159360, 3167741, 4229103, 1227493, 1401499, 1986134, 
    3211356, 4230788,
  1895025, 1230559, 2135147, 1092269, 1130181, 4241910, 775667, 16412, 
    3921076, 2327022 ;

 populationCity =
  1557980, 421014, 2945140, 13727, 3676953, 3581830, 1115203, 1791817, 
    4179906, 1642366,
  4675416, 2171007, 3434887, 601754, 2126773, 1258770, 2371912, 4374489, 
    1641720, 3782852,
  88046, 66073, 3842015, 1409696, 4172013, 3957536, 249425, 1870645, 3573016, 
    685060,
  2484579, 2686917, 3568779, 3711482, 3007543, 2813051, 1934855, 415058, 
    2900689, 4361222,
  4275846, 3935954, 3408511, 1785209, 4273344, 376844, 3481854, 2576121, 
    2398914, 3709248,
  548580, 309139, 4560466, 3814538, 2953378, 1664882, 1132587, 2293065, 
    2160044, 745202,
  766084, 3585058, 1325880, 2141219, 1534828, 1039834, 549413, 4602791, 
    2079739, 4615274,
  1137324, 3560275, 4458599, 932463, 2896950, 2476861, 2518382, 3190411, 
    933833, 247996,
  2918793, 4302224, 1358366, 742420, 1477456, 4014593, 1805771, 3781946, 
    2697613, 2341883,
  4097779, 729446, 3796200, 4444479, 2622899, 607349, 2755538, 1548797, 
    462074, 3898088 ;
}
